module accumulator(input clock,
						 input Ea,
						 input load_a,
						 inout logic [7:0] w_bus)
						 
endmodule
